/*
 * Copyright (c) 2020-2021, SERI Development Team
 *
 * SPDX-License-Identifier: Apache-2.0
 *
 * Change Logs:
 * Date           Author       Notes
 * 2022-01-26     Lyons        first version
 */

`include "pa_soc_param.v"

module M74HC154 (
    input  [3:0]                A,
    input  [1:0]                ENn,
           
    output [15:0]               Y
);

wire [15:0]                     TMP;

assign TMP[15:0] = {16{4'h0 == A[3:0]}} & 16'b1111_1111_1111_1110
                 | {16{4'h1 == A[3:0]}} & 16'b1111_1111_1111_1101
                 | {16{4'h2 == A[3:0]}} & 16'b1111_1111_1111_1011
                 | {16{4'h3 == A[3:0]}} & 16'b1111_1111_1111_0111
                 | {16{4'h4 == A[3:0]}} & 16'b1111_1111_1110_1111
                 | {16{4'h5 == A[3:0]}} & 16'b1111_1111_1101_1111
                 | {16{4'h6 == A[3:0]}} & 16'b1111_1111_1011_1111
                 | {16{4'h7 == A[3:0]}} & 16'b1111_1111_0111_1111
                 | {16{4'h8 == A[3:0]}} & 16'b1111_1110_1111_1111
                 | {16{4'h9 == A[3:0]}} & 16'b1111_1101_1111_1111
                 | {16{4'ha == A[3:0]}} & 16'b1111_1011_1111_1111
                 | {16{4'hb == A[3:0]}} & 16'b1111_0111_1111_1111
                 | {16{4'hc == A[3:0]}} & 16'b1110_1111_1111_1111
                 | {16{4'hd == A[3:0]}} & 16'b1101_1111_1111_1111
                 | {16{4'he == A[3:0]}} & 16'b1011_1111_1111_1111
                 | {16{4'hf == A[3:0]}} & 16'b0111_1111_1111_1111;

assign Y[15:0]   = (2'b00 == ENn[1:0]) ? TMP[15:0]
                                       : 16'b1111_1111_1111_1111;

endmodule